LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;


ENTITY DRIVER IS
	PORT(CTRL : IN STD_LOGIC;
		 D_OUT : OUT STD_LOGIC
	);
END ENTITY;

ARCHITECTURE BEHAVIORAL OF DRIVER IS

BEGIN

D_PROCESS: PROCESS(CTRL)
BEGIN
IF(CTRL = '1') THEN
	D_OUT <= 'Z';
	ELSE D_OUT <= '1';
END IF;
END PROCESS;

END ARCHITECTURE;
