LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY GENERICS_MUX IS
	GENERIC(INPUTS : INTEGER := 15; SIZE: INTEGER := 1); --N INPUT, N BIT
	PORT(INS : IN SIGNED((INPUTS*SIZE)-1 DOWNTO 0);
		 SEL : IN INTEGER;
		 OUT_MUX : OUT SIGNED(SIZE-1 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE BEH OF GENERICS_MUX IS
TYPE MATRIX IS ARRAY(0 TO INPUTS-1) OF SIGNED(SIZE - 1 DOWNTO 0);
SIGNAL MUX_IN : MATRIX;
BEGIN
  GEN : FOR I IN 0 TO INPUTS - 1 GENERATE
        MUX_IN(I) <= INS(((I + 1) * SIZE) - 1 DOWNTO (I * SIZE));
        END GENERATE;
    OUT_MUX <= MUX_IN(SEL);
END ARCHITECTURE;
