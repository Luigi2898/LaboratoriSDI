LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.all;

ENTITY DECODER IS
	PORT(W  : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 Y  : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 EN : IN STD_LOGIC	
	);
END ENTITY;

ARCHITECTURE BEHAVIOURAL OF DECODER IS

BEGIN

DEC : PROCESS(EN, W)
	 BEGIN
	     IF(EN = '1') THEN
	         CASE W IS
				 WHEN "0000" => Y <= STD_LOGIC_VECTOR(TO_UNSIGNED(0, 16));
				 WHEN "0001" => Y <= STD_LOGIC_VECTOR(TO_UNSIGNED(1, 16));
				 WHEN "0010" => Y <= STD_LOGIC_VECTOR(TO_UNSIGNED(2, 16));
				 WHEN "0011" => Y <= STD_LOGIC_VECTOR(TO_UNSIGNED(3, 16));
				 WHEN "0100" => Y <= STD_LOGIC_VECTOR(TO_UNSIGNED(4, 16));
				 WHEN "0101" => Y <= STD_LOGIC_VECTOR(TO_UNSIGNED(5, 16));
				 WHEN "0110" => Y <= STD_LOGIC_VECTOR(TO_UNSIGNED(6, 16));
				 WHEN "0111" => Y <= STD_LOGIC_VECTOR(TO_UNSIGNED(7, 16));
				 WHEN "1000" => Y <= STD_LOGIC_VECTOR(TO_UNSIGNED(8, 16));
				 WHEN "1001" => Y <= STD_LOGIC_VECTOR(TO_UNSIGNED(9, 16));
				 WHEN "1010" => Y <= STD_LOGIC_VECTOR(TO_UNSIGNED(10, 16));
				 WHEN "1011" => Y <= STD_LOGIC_VECTOR(TO_UNSIGNED(11, 16));
				 WHEN "1100" => Y <= STD_LOGIC_VECTOR(TO_UNSIGNED(12, 16));
				 WHEN "1101" => Y <= (OTHERS => 'Z');
				 WHEN "1110" => Y <= (OTHERS => 'Z');
				 WHEN "1111" => Y <= (OTHERS => 'Z');
				 WHEN OTHERS => Y <= (OTHERS => 'Z');
			END CASE;	 
	     END IF;
	 END PROCESS;
END ARCHITECTURE;