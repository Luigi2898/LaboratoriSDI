library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity multiplier is
  port (
  clock
  );
end entity;

architecture  of multiplier is

begin

end architecture;
