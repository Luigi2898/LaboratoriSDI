LIBRARY IEEE;
  USE IEEE.STD_LOGIC_1164.ALL;

ENTITY TB IS
END ENTITY;

ARCHITECTURE ARCH OF TB IS

  COMPONENT  RX IS
    PORT (
    CLK : IN STD_LOGIC;
    RST : IN STD_LOGIC;
    RX : IN STD_LOGIC;
    RD : IN STD_LOGIC;
    DATA : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    DAV : OUT STD_LOGIC
    );
  END COMPONENT;

  SIGNAL CLK : STD_LOGIC;
  SIGNAL RST : STD_LOGIC;
  SIGNAL RX1 : STD_LOGIC;
  SIGNAL RD : STD_LOGIC;
  SIGNAL DATA : STD_LOGIC_VECTOR(7 DOWNTO 0);
  SIGNAL DAV : STD_LOGIC;

BEGIN

  RIC : RX PORT MAP(CLK, RST, RX1, RD, DATA, DAV);

  CLOCK : PROCESS
  BEGIN

      CLK <= '0';
    WAIT FOR 20 NS;
      CLK <= '1';
    WAIT FOR 20 NS;
  END PROCESS;


  REST : PROCESS
  BEGIN
    RST <= '1';
    WAIT FOR 21 NS;
    RST <= '0';

  END PROCESS;

  RD <= '0';

  TRASMISSION : PROCESS
  BEGIN
    RX1 <= '1';
    WAIT FOR 50 NS;
    RX1 <= '0';
    WAIT FOR 104 US;
    RX1 <= '1';
    WAIT FOR 104 US;
    RX1 <= '0';
    WAIT FOR 104 US;
    RX1 <= '0';
    WAIT FOR 104 US;
    RX1 <= '1';
    WAIT FOR 104 US;
    RX1 <= '1';
    WAIT FOR 104 US;
    RX1 <= '0';
    WAIT FOR 104 US;
    RX1 <= '1';
    WAIT FOR 104 US;
    RX1 <= '0';
    WAIT FOR 104 US;
    RX1 <= '1';
  END PROCESS;
END ARCHITECTURE;
