LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY REG_N IS
GENERIC ( N : INTEGER := 8);
PORT(
		IN_REG : IN STD_LOGIC_VECTOR (N-1 DOWNTO 0);
		CLK, ENABLE, RST : IN STD_LOGIC;
		OUT_REG : OUT STD_LOGIC_VECTOR (N-1 DOWNTO 0)
	);
END REG_N;

ARCHITECTURE BEHAVIOUR OF REG_N IS
BEGIN

REG : PROCESS (CLK)
BEGIN
	IF (CLK'EVENT AND CLK = '1') THEN
		IF (RST = '0') THEN
			OUT_REG <= (OTHERS => '0');
		ELSIF (ENABLE = '1') THEN
			OUT_REG <= IN_REG;
		END IF;
	END IF;
END PROCESS;

END BEHAVIOUR;

