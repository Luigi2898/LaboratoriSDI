LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.all;

ENTITY MUX IS
	GENERIC(N : INTEGER := 47);
	PORT(IN_MUX, W_R, W_I : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		 OUT_MUX : OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		 SEL : IN STD_LOGIC_VECTOR(1 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE BEHAVIOURAL OF MUX IS

BEGIN

OUT_MUX <= IN_MUX WHEN SEL = "00" else
	            W_R WHEN SEL = "01" else
							W_I WHEN SEL = "10" else
							(others => 'Z');

END ARCHITECTURE;
