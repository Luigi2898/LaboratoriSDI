LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY UART IS

  PORT(
    DATA_IN  : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    TX_PIN   : OUT STD_LOGIC;
    TX_READY : OUT STD_LOGIC;
    WR       : IN STD_LOGIC;

    DATA_OUT : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    RX_PIN   : IN STD_LOGIC;
    RD       : IN STD_LOGIC;
    DAV      : OUT STD_LOGIC;

    CLOCK    : IN STD_LOGIC;
    RESETN   : IN STD_LOGIC
    );

END ENTITY;
 
ARCHITECTURE BEHAVIOURAL OF UART IS

  COMPONENT RX IS
    PORT (
      CLK  : IN STD_LOGIC;
      RST  : IN STD_LOGIC;
      RX   : IN STD_LOGIC;
      RD   : IN STD_LOGIC;
      DATA : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
      DAV  : OUT STD_LOGIC
    );
  END COMPONENT;

  COMPONENT TX IS
	 PORT(
     CLOCK       : IN STD_LOGIC;
		 RST         : IN STD_LOGIC;
		 DATA_IN     : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 TX          : OUT STD_LOGIC;
		 DATA_VALID  : IN STD_LOGIC;
		 TXREADY     : OUT STD_LOGIC
	 );
  END COMPONENT;

  BEGIN

    RECEIVER    : RX PORT MAP(CLOCK, RESETN, RX_PIN, RD, DATA_OUT, DAV);
    TRANSMITTER : TX PORT MAP(CLOCK, RESETN, DATA_IN, TX_PIN, WR, TX_READY);


END ARCHITECTURE;
