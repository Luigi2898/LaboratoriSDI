LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY FILTER_BLOCK IS
	port(CLK, RST : IN STD_LOGIC;
		 PDM : IN STD_LOGIC;
		 FILTERED : OUT SIGNED(13 DOWNTO 0)	
	);	

END ENTITY;

ARCHITECTURE BEH OF FILTER_BLOCK IS

COMPONENT FILTER IS
	PORT(PDM_IN, EN_CNT, CHIP_S : IN STD_LOGIC;
		 FILTERED : OUT SIGNED(13 DOWNTO 0);
		 CLK, RST : IN STD_LOGIC	
	);
END COMPONENT;

COMPONENT CU_FILTER IS
	PORT(CLK, RST : IN STD_LOGIC;
		 EN_CNT, CHIP_S, FILT_RST : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL EN_CNT, CHIP_S, FILT_RST : STD_LOGIC;

BEGIN
FIL: FILTER PORT MAP(PDM, EN_CNT, CHIP_S, FILTERED, CLK, FILT_RST);
CU : CU_FILTER PORT MAP(CLK, RST, EN_CNT, CHIP_S, FILT_RST);



END ARCHITECTURE;