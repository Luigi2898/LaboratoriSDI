LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY PL_REG_N IS
GENERIC ( N_BIT : INTEGER := 8);
PORT(
		IN_REG : IN STD_LOGIC_VECTOR (N_BIT-1 DOWNTO 0);
		CLK, ENABLE, CLR : IN STD_LOGIC;
		OUT_REG : OUT STD_LOGIC_VECTOR (N_BIT-1 DOWNTO 0)
	);
END PL_REG_N;

ARCHITECTURE BEHAVIOUR OF PL_REG_N IS
BEGIN

TRANSFER_PROCESS : PROCESS (CLK)
BEGIN
	IF (CLK'EVENT AND CLK = '1') THEN
		IF (CLR = '0') THEN
			OUT_REG <= (OTHERS => '0');
		ELSIF (ENABLE = '1') THEN
			OUT_REG <= IN_REG;
		END IF;
	END IF;
END PROCESS;

END BEHAVIOUR;

