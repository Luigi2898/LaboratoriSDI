LIBRARY IEEE;
  USE IEEE.STD_LOGIC_1164.ALL;

ENTITY  RX IS
  PORT (
  CLK : IN STD_LOGIC;
  RST : IN STD_LOGIC;
  RX : IN STD_LOGIC;
  RD : IN STD_LOGIC;
  DATA : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
  DAV : OUT STD_LOGIC
  );
END ENTITY;

ARCHITECTURE BEHAVIOURAL OF RX IS
  COMPONENT CU_RX IS
  	PORT(CLOCK          : IN STD_LOGIC;
           RST            : IN STD_LOGIC;
  		 S_BIT          : IN STD_LOGIC;
  		 DATA_VALID     : OUT STD_LOGIC;
  		 DP_RST         : OUT STD_LOGIC;
  		 RD             : IN STD_LOGIC;
  		 BAUD_EN        : OUT STD_LOGIC;
  		 BAUD_END       : IN  STD_LOGIC;
  		 FRAME_EN       : OUT STD_LOGIC;
  		 FRAME_END      : IN STD_LOGIC;
       FRAME_RST : OUT STD_LOGIC;
  	     ENABLE_INPUT   : OUT STD_LOGIC;
  		 ENABLE_OUTPUT  : OUT STD_LOGIC
  	);
  END COMPONENT;

  COMPONENT DP IS
    PORT (
    RX : IN STD_LOGIC;
    RST :  IN STD_LOGIC;
    CLOCK : IN STD_LOGIC;
    ENINPUT : IN STD_LOGIC;
    STARTBIT : OUT STD_LOGIC;
    EN_OUT_REG : IN STD_LOGIC;
    DATAOUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    BAUD_EN : IN STD_LOGIC;
    BAUD_END : OUT STD_LOGIC;
    FRAME_EN : IN STD_LOGIC;
    FRAME_END : OUT STD_LOGIC;
    FRAME_RST : IN STD_LOGIC
    );
  END COMPONENT;

  SIGNAL ENINPUT : STD_LOGIC;
  SIGNAL STARTBIT : STD_LOGIC;
  SIGNAL EN_OUT_REG : STD_LOGIC;
  SIGNAL  BAUD_EN : STD_LOGIC;
  SIGNAL BAUD_END : STD_LOGIC;
  SIGNAL  FRAME_EN : STD_LOGIC;
  SIGNAL FRAME_END : STD_LOGIC;
  SIGNAL DP_RESET : STD_LOGIC;
  SIGNAL FRAME_RST : STD_LOGIC;

BEGIN

  DADATAPATH : DP PORT MAP(RX, DP_RESET, CLK, ENINPUT, STARTBIT, EN_OUT_REG, DATA, BAUD_EN, BAUD_END, FRAME_EN, FRAME_END, FRAME_RST);
  CONTROL_UNIT : CU_RX PORT MAP(CLK, RST, STARTBIT, DAV, DP_RESET, RD, BAUD_EN, BAUD_END, FRAME_EN, FRAME_END, FRAME_RST, ENINPUT, EN_OUT_REG);

END ARCHITECTURE;
