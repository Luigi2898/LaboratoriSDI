LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY TX IS
	PORT(CLOCK       : IN STD_LOGIC;
		 RST         : IN STD_LOGIC;
		 DATA_IN     : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 TX          : OUT STD_LOGIC;
		 DATA_VALID  : IN STD_LOGIC;
		 TXREADY     : OUT STD_LOGIC	
	);
END ENTITY;


ARCHITECTURE STRUCT OF TX IS

COMPONENT DP_TX IS
	PORT(CLOCK     : IN STD_LOGIC;
		 DATA_IN   : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 BAUD_END  : OUT STD_LOGIC;
		 SHIFT_END : OUT STD_LOGIC;
		 SH_OUT    : OUT STD_LOGIC;
		 DP_RST    : IN STD_LOGIC;
		 BAUD_CNT  : IN STD_LOGIC;
		 SHIFT_CNT : IN STD_LOGIC;
		 SHIFT_EN  : IN STD_LOGIC;
		 LOAD_EN   : IN STD_LOGIC;
		 READ_EN   : IN STD_LOGIC	
	);
END COMPONENT;

COMPONENT CU IS
  PORT (
    CLOCK      : IN STD_LOGIC;
    RST        : IN STD_LOGIC;
    BAUD_END   : IN STD_LOGIC;
    SHIFT_END  : IN STD_LOGIC;
    DATA_VALID : IN STD_LOGIC;
    DP_RST     : OUT STD_LOGIC;
    BAUD_CNT   : OUT STD_LOGIC;
    SHIFT_CNT  : OUT STD_LOGIC;
    SHIFT_EN   : OUT STD_LOGIC;
    LOAD_EN    : OUT STD_LOGIC;
    READ_EN    : OUT STD_LOGIC;
    TXREADY    : OUT STD_LOGIC
  );
END COMPONENT;

SIGNAL BAUD_END, SHIFT_END, SH_OUT, BAUD_CNT, SHIFT_CNT, SHIFT_EN, LOAD_EN, RD_EN, DP_RST : STD_LOGIC;

BEGIN
DP : DP_TX PORT MAP(CLOCK, DATA_IN, BAUD_END, SHIFT_END, TX, DP_RST, BAUD_CNT, SHIFT_CNT, SHIFT_EN, LOAD_EN, RD_EN);

CONTROL : CU PORT MAP(CLOCK, RST, BAUD_END, SHIFT_END, DATA_VALID, DP_RST, BAUD_CNT, SHIFT_CNT, SHIFT_EN, LOAD_EN, RD_EN, TXREADY);

END ARCHITECTURE;
