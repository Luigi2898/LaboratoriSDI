LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY CU_FILTER IS
	PORT(CLK, RST : IN STD_LOGIC;
		 EN_CNT, CHIP_S, FILT_RST : OUT STD_LOGIC
	);
END ENTITY;

ARCHITECTURE BEH OF CU_FILTER IS

TYPE STATE_TYPE IS (RST_S, IDLE);
SIGNAL STATE : STATE_TYPE;

BEGIN
FSM : PROCESS(CLK, RST)
BEGIN
IF(RST = '0') THEN
	STATE <= RST_S;
	ELSIF(CLK'EVENT AND CLK = '1') THEN
		CASE(STATE) IS
			WHEN RST_S => STATE <= IDLE;
			WHEN IDLE => STATE <= IDLE;
			WHEN OTHERS => STATE <= RST_S;
		END CASE;
END IF;
END PROCESS;	

OUTPUT : PROCESS(STATE)
BEGIN
FILT_RST <= '1';
EN_CNT <= '0';
CHIP_S <= '0';
CASE (STATE) IS
	WHEN RST_S => 
		 FILT_RST <= '0';
	WHEN IDLE =>
		 EN_CNT <= '1';
	     CHIP_S <= '1';
END CASE;
END PROCESS;

END ARCHITECTURE;
