LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;


ENTITY CU_FRONT_END IS
	PORT(CLK_10N : IN STD_LOGIC;
	     CLK_MIC  : IN STD_LOGIC;
		 RST_CU     : IN STD_LOGIC;
		 RST_CNT1 : OUT STD_LOGIC;
		 RST_CNT2  : OUT STD_LOGIC;
		 TC_HIGH : IN STD_LOGIC;
		 TC_HIGN_NEG : IN STD_LOGIC;
		 FF_IN : OUT STD_LOGIC;
		 EN_FF1 : OUT STD_LOGIC;
		 RST_FF1: OUT STD_LOGIC;
		 FF_IN_NEG : OUT STD_LOGIC;
		 EN_FF2  : OUT STD_LOGIC;
		 RST_FF2 : OUT STD_LOGIC
	);
END ENTITY;

ARCHITECTURE BEH OF CU_FRONT_END IS

TYPE STATE_HIGH IS (IDLE1, COUNT1, SET1, RESET_FF1);
TYPE STATE_LOW IS (IDLE2, COUNT2, SET2, RESET_FF2);
SIGNAL STATE1 : STATE_HIGH;
SIGNAL STATE2 : STATE_LOW;
SIGNAL CLK_MIC_N : STD_LOGIC;

BEGIN
CLK_MIC_N <= NOT(CLK_MIC);

STATE_P1: PROCESS(CLK_10N, CLK_MIC, RST_CU)
BEGIN
IF(RST_CU = '0') THEN
  STATE1 <= IDLE1;
  ELSIF(CLK_10N = '1' AND CLK_10N'EVENT) THEN
     CASE STATE1 IS
	 WHEN IDLE1 => IF(CLK_MIC = '1') THEN
				   STATE1 <= COUNT1;
				   ELSE STATE1 <= IDLE1;
				   END IF;
	 WHEN COUNT1 => IF(TC_HIGH = '1') THEN
                   STATE1 <= SET1;
				   ELSE STATE1 <= COUNT1;
				   END IF;
     WHEN SET1 => STATE1 <= RESET_FF1;
	 WHEN RESET_FF1 => STATE1 <= IDLE1;
     WHEN OTHERS => STATE1 <= IDLE1;	 
	 END CASE;
END IF;
END PROCESS;


STATE_P2: PROCESS(CLK_10N, CLK_MIC_N, RST_CU)
BEGIN
IF(RST_CU = '0') THEN
  STATE2 <= IDLE2;
  ELSIF(CLK_10N = '1' AND CLK_10N'EVENT) THEN
     CASE STATE2 IS
	 WHEN IDLE2 => IF(CLK_MIC_N = '1') THEN
				   STATE2 <= COUNT2;
				   ELSE STATE2 <= IDLE2;
				   END IF;
	 WHEN COUNT2 => IF(TC_HIGN_NEG = '1') THEN
                   STATE2 <= SET2;
				   ELSE STATE2 <= COUNT2;
				   END IF;
     WHEN SET2 => STATE2 <= RESET_FF2;
	 WHEN RESET_FF2 => STATE2 <= IDLE2;
     WHEN OTHERS => STATE2 <= IDLE2;	 
	 END CASE;
END IF;
END PROCESS;


OUT_P1 : PROCESS(STATE1)
BEGIN
FF_IN <= '0';
EN_FF1 <= '0';
RST_FF1 <= '0';
RST_CNT1 <= '1';
CASE STATE1 IS
     WHEN IDLE1 => 
	 RST_FF1 <= '1'; 
     RST_CNT1 <= '0';
	 WHEN COUNT1 =>
	 EN_FF1 <= '1';
	 WHEN SET1 =>
	 FF_IN <= '1';
	 WHEN RESET_FF1 =>
	 
END CASE;
END PROCESS;

OUT_P2 : PROCESS(STATE2)
BEGIN
FF_IN_NEG <= '0';
EN_FF2 <= '0';
RST_FF2 <= '0';
RST_CNT2 <= '1';

CASE STATE2 IS
     WHEN IDLE2 => 
	 RST_FF2 <= '1'; 
     RST_CNT2 <= '0';
	 WHEN COUNT2 =>
	 EN_FF2 <= '1';
	 WHEN SET2 =>
	 FF_IN_NEG <= '1';
	 WHEN RESET_FF2 =>
	 
END CASE;
END PROCESS;





END ARCHITECTURE;
