LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY DP_DELAY IS
	PORT(CLK           : IN STD_LOGIC;
		 RST_DP        : IN STD_LOGIC;
		 EN_CNT_DELAY  : IN STD_LOGIC;
		 RST_CNT_DELAY : IN STD_LOGIC;
		 EN_FIRST      : IN STD_LOGIC;
	   EN_SECOND     : IN STD_LOGIC;
	   DELAY_END     : OUT STD_LOGIC;
		 DELAY_OUT     : BUFFER SIGNED(9 DOWNTO 0); --AGGIUNGERE BIT
     MSB           : OUT STD_LOGIC;
		 EN_DELAY_OUT  : IN STD_LOGIC;
		 SUB           : IN STD_LOGIC
	);
END ENTITY;

ARCHITECTURE BEH OF DP_DELAY IS

COMPONENT N_COUNTER IS
		GENERIC(N : INTEGER:= 6; MODULE : INTEGER := 42);
		PORT(CLK : IN STD_LOGIC;
			 EN  : IN STD_LOGIC;
			 RST : IN STD_LOGIC;
			 CNT_END : OUT STD_LOGIC;
			 CNT_OUT : BUFFER UNSIGNED(N-1 DOWNTO 0)
		);
END COMPONENT;

COMPONENT REG IS
	GENERIC(N : INTEGER := 8);
	PORT(REG_IN : IN signed(N-1 DOWNTO 0);
		 REG_OUT : OUT signed(N-1 DOWNTO 0);
		 CLK, RST, LOAD : IN STD_LOGIC
	);
END COMPONENT;

COMPONENT ADD_SUB IS
	GENERIC(N_AS : INTEGER := 20);
	PORT(IN_AS_1, IN_AS_2 : IN SIGNED(N_AS-1 DOWNTO 0);
		 AS_OUT : OUT SIGNED(N_AS-1 DOWNTO 0);
		 PDM: IN std_logic
	);
END COMPONENT;

SIGNAL CAPTURE : UNSIGNED(9 DOWNTO 0);
SIGNAL DELAY_AS  : SIGNED(9 DOWNTO 0);
SIGNAL DELAY1, DELAY2 : SIGNED(9 DOWNTO 0);
BEGIN

COUNT_DELAY: N_COUNTER GENERIC MAP(N => 10, MODULE => 1024) PORT MAP(CLK, EN_CNT_DELAY, RST_CNT_DELAY, DELAY_END, CAPTURE);

FIRST  : REG GENERIC MAP(N => 10) PORT MAP(SIGNED(CAPTURE), DELAY1, CLK, RST_DP, EN_FIRST);
SECOND : REG GENERIC MAP(N => 10) PORT MAP(SIGNED(CAPTURE), DELAY2, CLK, RST_DP, EN_SECOND);

AS_DELAY : ADD_SUB GENERIC MAP(N_AS => 10) PORT MAP(DELAY1, DELAY2, DELAY_AS, SUB);

out_delay : REG GENERIC MAP(N => 10) PORT MAP(DELAY_AS, DELAY_OUT, CLK, RST_DP, EN_DELAY_OUT);
MSB <= DELAY_OUT(9);


END ARCHITECTURE;
