library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity  is
  port (
  clock
  );
end entity;

architecture arch of  is

begin

end architecture;
