LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY VOTER IS
  PORT (

  IN1 : IN STD_LOGIC;
  IN2 : IN STD_LOGIC;
  IN3 : IN STD_LOGIC;
  WINNER : OUT STD_LOGIC

  );
END ENTITY;

ARCHITECTURE BEHAVIOURAL OF  VOTER IS

BEGIN

  WINNER <= (IN1 AND IN2) OR (IN1 AND IN3) OR (IN2 AND IN3);

END ARCHITECTURE;
