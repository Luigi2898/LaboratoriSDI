LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY ADD_SUB IS
	GENERIC(N_AS : INTEGER := 20);
	PORT(IN_AS_1, IN_AS_2 : IN SIGNED(N_AS-1 DOWNTO 0);
		 AS_OUT : OUT SIGNED(N_AS-1 DOWNTO 0);
		 PDM: IN std_logic
	);
END ENTITY;

ARCHITECTURE BEH OF ADD_SUB IS

SIGNAL IN1_NEG, IN2_NEG : SIGNED(N_AS-1 DOWNTO 0);	

BEGIN --ARCHITECTURE

PROCESS(IN_AS_1, IN_AS_2, PDM)
BEGIN
	IF(PDM = '1') THEN
	 AS_OUT <= IN_AS_1 + IN_AS_2;
	 ELSE AS_OUT <= IN_AS_1 - IN_AS_2;
    END IF; 
END PROCESS;


END ARCHITECTURE;