LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY FILTER IS
	PORT(PDM_IN, EN_CNT, CHIP_S : IN STD_LOGIC;
		 FILTERED : OUT SIGNED(13 DOWNTO 0);
		 CLK, RST : IN STD_LOGIC	
	);
END ENTITY;


ARCHITECTURE BEH OF FILTER IS

COMPONENT ROM IS
  PORT (
	CLK, CHIP_S : IN STD_LOGIC;
    ADDRESS : IN UNSIGNED(5 DOWNTO 0); 
    DATA    : OUT SIGNED(13 DOWNTO 0)
  );
END COMPONENT;

COMPONENT ADD_SUB IS
	GENERIC(N_AS : INTEGER := 14);
	PORT(IN_AS_1, IN_AS_2 : IN SIGNED(N_AS-1 DOWNTO 0);
		 AS_OUT : OUT SIGNED(N_AS-1 DOWNTO 0);
		 PDM: IN STD_LOGIC
	);

END COMPONENT;

COMPONENT REG IS
	PORT(REG_IN : IN STD_LOGIC;
		 REG_OUT : OUT STD_LOGIC;
		 CLK, RST : IN STD_LOGIC	
	);
END COMPONENT;

COMPONENT ACC IS 
	GENERIC(N_ACC : INTEGER := 14);
	PORT(ACC_IN : IN SIGNED(N_ACC-1 DOWNTO 0);
		 ACC_OUT : OUT SIGNED(N_ACC-1 DOWNTO 0);
		 CLK, RST: IN STD_LOGIC	
	);
END COMPONENT;



COMPONENT N_COUNTER IS
		GENERIC(N : INTEGER:= 6);
		PORT(CLK : IN STD_LOGIC;
			 EN  : IN STD_LOGIC;
			 RST : IN STD_LOGIC;
			 CNT_END : OUT STD_LOGIC;
			 CNT_OUT : BUFFER UNSIGNED(N-1 DOWNTO 0)		
		);
END COMPONENT;

SIGNAL CNT_END, REG_OUT: STD_LOGIC;
SIGNAL CNT_OUT: UNSIGNED(5 DOWNTO 0);
SIGNAL COEFF, ACC_OUT, AS_OUT : SIGNED(13 DOWNTO 0);
BEGIN

R1: REG PORT MAP(PDM_IN, REG_OUT, CLK, RST);
AS : ADD_SUB GENERIC MAP(N_AS => 14) PORT MAP(COEFF, ACC_OUT, AS_OUT, REG_OUT);
ACC1 : ACC GENERIC MAP(N_ACC => 14) PORT MAP(AS_OUT, ACC_OUT, CLK, RST);
CNT : N_COUNTER GENERIC MAP(N => 6) PORT MAP(CLK, EN_CNT, RST, CNT_END, CNT_OUT);
MEM : ROM PORT MAP(CLK, CHIP_S, CNT_OUT, COEFF);

FILTERED <= ACC_OUT;

END ARCHITECTURE;