LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY UARTQP IS

	PORT(
		SW : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		GPIO_0 : OUT STD_LOGIC_VECTOR(35 DOWNTO 0);
		KEY : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		LEDR : OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
		CLOCK_50 : IN STD_LOGIC
	);

END ENTITY;

ARCHITECTURE BEH OF UARTQP IS

  COMPONENT UART IS

    PORT(
      DATA_IN  : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      TX_PIN       : OUT STD_LOGIC;
      TX_READY : OUT STD_LOGIC;
      WR       : IN STD_LOGIC;

      DATA_OUT : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      RX_PIN       : IN STD_LOGIC;
      RD       : IN STD_LOGIC;
      DAV      : OUT STD_LOGIC;

      CLOCK    : IN STD_LOGIC;
      RESETN   : IN STD_LOGIC
    );

  END COMPONENT;


COMPONENT PLL IS
	PORT (
		REFCLK   : IN  STD_LOGIC := '0'; --  REFCLK.CLK
		RST      : IN  STD_LOGIC := '0'; --   RESET.RESET
		OUTCLK_0 : OUT STD_LOGIC;        -- OUTCLK0.CLK
		LOCKED   : OUT STD_LOGIC         --  LOCKED.EXPORT
	);
END COMPONENT PLL;

COMPONENT RISINGEDGE_DFLIPFLOP IS
   PORT(
      Q : OUT STD_LOGIC;
      CLK :IN STD_LOGIC;
      D :IN  STD_LOGIC
   );
END COMPONENT RISINGEDGE_DFLIPFLOP;

  SIGNAL TX, RD                    : STD_LOGIC;
  SIGNAL TX_READY  : STD_LOGIC;

  SIGNAL WR : STD_LOGIC ;

  SIGNAL D, D1 : STD_LOGIC;
  SIGNAL Q, Q1 : STD_LOGIC;

  SIGNAL CLOCK, OUTCLK_0, LOCKED  : STD_LOGIC;
  SIGNAL RESETN1, RESETN2      : STD_LOGIC;

BEGIN

  UART1 : UART PORT MAP (SW(7 DOWNTO 0), TX, GPIO_0(8), WR, LEDR(7 DOWNTO 0), TX, RD, GPIO_0(16), OUTCLK_0, KEY(2));
  GPIO_0(2) <= OUTCLK_0;
  GPIO_0(34) <= WR;
  GPIO_0(22) <= TX;
  GPIO_0(10) <= RD;
  --GPIO_0(10) <= KEY(2);

  PLLLL : PLL PORT MAP(CLOCK_50, NOT(KEY(2)), OUTCLK_0, LOCKED);

  FF : RISINGEDGE_DFLIPFLOP PORT MAP(Q, OUTCLK_0, D);
  FF1 : RISINGEDGE_DFLIPFLOP PORT MAP(Q1, OUTCLK_0, D1);

  KEYPROPC1 : PROCESS(KEY(0), OUTCLK_0)

  BEGIN
	IF(KEY(0)'EVENT AND KEY(0) = '0') THEN
		IF (OUTCLK_0 = '1') THEN
			WR <= '1';
			D <= '1';
		END IF;
	END IF;
	IF(OUTCLK_0 = '1' AND Q = '1') THEN
		WR <= '0';
		D <= '0';
	END IF;
  END PROCESS;

  KEYPROPC2 : PROCESS(KEY(1), OUTCLK_0)

  BEGIN
	IF(KEY(1)'EVENT AND KEY(1) = '0') THEN
		IF (OUTCLK_0 = '1') THEN
			RD <= '1';
			D1 <= '1';
		END IF;
	END IF;
	IF(OUTCLK_0 = '1' AND Q1 = '1') THEN
		RD <= '0';
		D1 <= '0';
	END IF;
  END PROCESS;



END ARCHITECTURE;
