LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY REG IS
	PORT(REG_IN : IN STD_LOGIC;
		 REG_OUT : OUT STD_LOGIC;
		 CLK, RST, LOAD : IN STD_LOGIC	
	);
END ENTITY;

ARCHITECTURE BEH OF REG IS

BEGIN
REGPROC: PROCESS(CLK)
BEGIN
IF(RST = '0') THEN
	REG_OUT <= '0';
     ELSIF(CLK'EVENT AND CLK = '1') THEN
		 IF(LOAD = '1') THEN
		 REG_OUT <= REG_IN;
		 END IF;
END IF;

END PROCESS;

END ARCHITECTURE;