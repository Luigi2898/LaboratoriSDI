LIBRARY IEEE;
  USE IEEE.STD_LOGIC_1164.ALL;
  USE IEEE.NUMERIC_STD.ALL;

--DATAPATH RX

ENTITY DP IS
  PORT (RX         : IN  STD_LOGIC;
        RST        : IN  STD_LOGIC;
        CLOCK      : IN  STD_LOGIC;
        ENINPUT    : IN  STD_LOGIC;
        STARTBIT   : OUT STD_LOGIC;
        EN_OUT_REG : IN  STD_LOGIC;
        DATAOUT    : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
        BAUD_EN    : IN  STD_LOGIC;
        BAUD_END   : OUT STD_LOGIC;
        FRAME_EN   : IN  STD_LOGIC;
        FRAME_END  : OUT STD_LOGIC;
        FRAME_RST  : IN  STD_LOGIC
  );
END ENTITY;

ARCHITECTURE BEHAVIOURAL OF DP IS

  COMPONENT N_COUNTER IS
  		GENERIC(N      : INTEGER:= 12;
              MODULE : INTEGER:= 2604);
  		PORT(CLK     : IN STD_LOGIC;
  			   EN      : IN STD_LOGIC;
  			   RST     : IN STD_LOGIC;
  			   CNT_END : OUT STD_LOGIC;
  			   CNT_OUT : BUFFER UNSIGNED(N-1 DOWNTO 0)
  		);
  END COMPONENT;

  COMPONENT SERIAL2PARALLEL IS
  GENERIC(N : INTEGER);
  	PORT(CLK        : IN STD_LOGIC;
  		   RST        : IN STD_LOGIC;
  		   EN         : IN STD_LOGIC;
  		   SERIAL_D   : IN STD_LOGIC;
  		   PARALLEL_D : BUFFER STD_LOGIC_VECTOR(N-1 DOWNTO 0)
  	);
  END COMPONENT;

  COMPONENT STARTBITFINDER IS
    PORT (
      FRAME : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      STARTBIT : OUT STD_LOGIC
    );
  END COMPONENT;

  COMPONENT VOTER IS
    PORT (
    IN1 : IN STD_LOGIC;
    IN2 : IN STD_LOGIC;
    IN3 : IN STD_LOGIC;
    WINNER : OUT STD_LOGIC
    );
  END COMPONENT;

  SIGNAL BAUD_COUNT_OUT  : UNSIGNED(11 DOWNTO 0);
  SIGNAL FRAME_COUNT_OUT : UNSIGNED(2 DOWNTO 0);
  SIGNAL TO_LOGIC        : STD_LOGIC_VECTOR(7 DOWNTO 0);
  SIGNAL VOTE            : STD_LOGIC;
  SIGNAL IN1, IN2, IN3   : STD_LOGIC;

BEGIN

  BAUD_COUNTER  : N_COUNTER       GENERIC MAP(12, 2604)
                                  PORT MAP(CLOCK, BAUD_EN, RST, BAUD_END, BAUD_COUNT_OUT);
  FRAME_COUNTER : N_COUNTER       GENERIC MAP(3, 7)
                                  PORT MAP(CLOCK, FRAME_EN, FRAME_RST, FRAME_END, FRAME_COUNT_OUT);
  INPUT_REG     : SERIAL2PARALLEL GENERIC MAP(8)
                                  PORT MAP(CLOCK, RST, ENINPUT, RX, TO_LOGIC);
  OUTPUT_REG    : SERIAL2PARALLEL GENERIC MAP(8)
                                  PORT MAP(CLOCK, RST, EN_OUT_REG , VOTE , DATAOUT);
  VOTATORE      : VOTER           PORT MAP(TO_LOGIC(3), TO_LOGIC(4), TO_LOGIC(5), VOTE);

  S_BIT_F       : STARTBITFINDER  PORT MAP(TO_LOGIC, STARTBIT);

END ARCHITECTURE;
