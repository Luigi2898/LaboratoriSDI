LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY REG IS
	GENERIC(N : INTEGER := 8);
	PORT(REG_IN : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		 REG_OUT : OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		 CLK, RST, LOAD : IN STD_LOGIC	
	);
END ENTITY;

ARCHITECTURE BEH OF REG IS

BEGIN
REGPROC: PROCESS(CLK, RST)
BEGIN
IF(RST = '0') THEN
	REG_OUT <= (OTHERS => '0');
     ELSIF(CLK'EVENT AND CLK = '1') THEN
		 IF(LOAD = '1') THEN
		 REG_OUT <= REG_IN;
		 END IF;
END IF;

END PROCESS;

END ARCHITECTURE;