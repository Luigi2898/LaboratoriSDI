LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;


ENTITY POLYPHASE_FIR IS
	GENERIC(INITFILE : STRING := "POLYPHASE.TXT");
	PORT(CLK      : IN STD_LOGIC;
	     RST      : IN STD_LOGIC;
	     DOWNS_IN : IN STD_LOGIC;
	     M_DIV_END: IN STD_LOGIC;
		 DAV      : OUT STD_LOGIC;
		 FIR_OUT  : BUFFER SIGNED(23 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE BEH OF POLYPHASE_FIR IS 

COMPONENT FIR IS
	GENERIC(INITFILE : STRING := "POLYPHASE.TXT");
	PORT(CLK         : IN STD_LOGIC; 
	     RST_FIR     : IN STD_LOGIC;
		 RST_CNT_FIR : IN STD_LOGIC;
	     EN_CNT_FIR  : IN STD_LOGIC; 		 
		 DOWNS_IN    : IN STD_LOGIC;
		 CNT_END_POLY: OUT STD_LOGIC; 	
		 OUT_MUX     : OUT STD_LOGIC_VECTOR(0 DOWNTO 0); 
		 PDM_AS      : IN STD_LOGIC;
		 EN_ACC      : IN STD_LOGIC;
		 RST_ACC     : IN STD_LOGIC;
		 LOAD_EN     : IN STD_LOGIC; 
		 SHIFT_EN    : IN STD_LOGIC; 
		 FIR_OUT     : BUFFER SIGNED(23 DOWNTO 0) 
	);
END COMPONENT;

COMPONENT CU_POLYPHASE IS 
	PORT(CLK         : IN STD_LOGIC;
         RST         : IN STD_LOGIC;
		 RST_FIR     : OUT STD_LOGIC;
		 RST_CNT_FIR : OUT STD_LOGIC;
		 EN_CNT_FIR  : OUT STD_LOGIC;
		 CNT_END_POLY: IN STD_LOGIC;
		 OUT_MUX     : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
		 PDM_AS	     : OUT STD_LOGIC;
		 EN_ACC      : OUT STD_LOGIC;
		 RST_ACC     : OUT STD_LOGIC;
		 LOAD_EN     : OUT STD_LOGIC;
		 DAV	     : OUT STD_LOGIC;
		 SHIFT_EN    : OUT STD_LOGIC; 
		 M_DIV_END   : IN STD_LOGIC		 	
	);
END COMPONENT;

SIGNAL EN_CNT_FIR, CNT_END_POLY, PDM_AS, EN_ACC, RST_ACC, LOAD_EN, RST_FIR, RST_CNT_FIR, SHIFT_EN : STD_LOGIC;
SIGNAL OUT_MUX : STD_LOGIC_VECTOR(0 DOWNTO 0);

BEGIN
FIR0 : FIR GENERIC MAP(INITFILE => INITFILE) PORT MAP(CLK, RST_FIR, RST_CNT_FIR, EN_CNT_FIR, DOWNS_IN, CNT_END_POLY, 
													  OUT_MUX, PDM_AS, EN_ACC, RST_ACC, LOAD_EN, SHIFT_EN, FIR_OUT);

CU : CU_POLYPHASE PORT MAP(CLK, RST, RST_FIR, RST_CNT_FIR, EN_CNT_FIR, CNT_END_POLY, 
                           OUT_MUX, PDM_AS, EN_ACC, RST_ACC, LOAD_EN, DAV, SHIFT_EN, M_DIV_END); 

END ARCHITECTURE;