LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY FILTER IS
	PORT(CLK           : IN STD_LOGIC;
         RST_ALL       : IN STD_LOGIC;
	     PDM_IN        : IN STD_LOGIC;
		 LOAD          : IN STD_LOGIC;
		 M_EN          : IN STD_LOGIC;
		 DAV_OUT       : OUT STD_LOGIC_VECTOR(7 DOWNTO 0); --MANDARE ALLA CU
		 DAV_IN        : IN STD_LOGIC; --DALLA CU PER SOMMARE TUTTO
		 POLY_VALID    : IN STD_LOGIC;
		 EN_CNT_ADD    : IN STD_LOGIC;
		 RST_ACC       : IN STD_LOGIC;
		 EN_ACC        : IN STD_LOGIC;
		 RST_M_DIV     : IN STD_LOGIC;
		 M_DIV_END_IN  : IN STD_LOGIC; --DALLA CU
		 M_DIV_END_OUT : OUT STD_LOGIC; --ALLA CU
		 CNT_END       : OUT STD_LOGIC; --ALLA CU
	     FILTER_OUT    : BUFFER SIGNED(27 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE BEH OF FILTER IS

COMPONENT POLYPHASE_FIR IS
	GENERIC(INITFILE : STRING := "POLYPHASE.TXT");
	PORT(CLK         :IN STD_LOGIC;
	     RST         : IN STD_LOGIC;
	     DOWNS_IN    : IN STD_LOGIC;
	     M_DIV_END   : IN STD_LOGIC;
		 DAV         : OUT STD_LOGIC;
		 POLY_VALID  : IN STD_LOGIC;
		 FIR_OUT     : BUFFER SIGNED(27 DOWNTO 0)
	);
END COMPONENT;

COMPONENT N_COUNTER IS
    GENERIC(N : INTEGER:= 6; MODULE : INTEGER := 42);
	PORT(CLK : IN STD_LOGIC;
		 EN  : IN STD_LOGIC;
		 RST : IN STD_LOGIC;
		 CNT_END : OUT STD_LOGIC;
		 CNT_OUT : BUFFER UNSIGNED(N-1 DOWNTO 0)		
	);
END COMPONENT;

COMPONENT FF IS
	PORT(FF_IN : IN STD_LOGIC;
		 FF_OUT : OUT STD_LOGIC;
		 CLK, RST, LOAD : IN STD_LOGIC	
	);
END COMPONENT;

COMPONENT ADD_SUB IS
	GENERIC(N_AS : INTEGER := 20);
	PORT(IN_AS_1, IN_AS_2 : IN SIGNED(N_AS-1 DOWNTO 0);
		 AS_OUT : OUT SIGNED(N_AS-1 DOWNTO 0);
		 PDM: IN std_logic
	);
END COMPONENT;

COMPONENT ACC IS 
	GENERIC(N_ACC : INTEGER := 14);
	PORT(ACC_IN : IN SIGNED(N_ACC-1 DOWNTO 0);
		 ACC_OUT : OUT SIGNED(N_ACC-1 DOWNTO 0);
		 CLK, RST, EN_ACC: IN STD_LOGIC	
	);
END COMPONENT;


COMPONENT GENERICS_MUX IS
	GENERIC(INPUTS : INTEGER := 15; SIZE: INTEGER := 1); --N INPUT, N BIT 
	PORT(INS : IN STD_LOGIC_VECTOR((INPUTS*SIZE)-1 DOWNTO 0);
		 SEL : IN INTEGER;
		 OUT_MUX : OUT STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0)
	);
END COMPONENT;


SIGNAL M_OUT: UNSIGNED(2 DOWNTO 0);
SIGNAL REG_OUT: STD_LOGIC_VECTOR(6 DOWNTO 0); --OUT Z_REG  
SIGNAL AS_OUT : SIGNED(27 DOWNTO 0);
SIGNAL P_OUT0,P_OUT1,P_OUT2,P_OUT3,P_OUT4, P_OUT5, P_OUT6, P_OUT7: SIGNED(27 DOWNTO 0);
SIGNAL DAV0, DAV1, DAV2, DAV3, DAV4, DAV5, DAV6, DAV7 : STD_LOGIC;
SIGNAL P_IN_MUX : SIGNED(223 DOWNTO 0);
SIGNAL P_OUT_MUX: STD_LOGIC_VECTOR(27 DOWNTO 0);
SIGNAL CNT_OUT: UNSIGNED(2 DOWNTO 0);
BEGIN

M_DIVIDER : N_COUNTER GENERIC MAP(N => 3, MODULE => 8) PORT MAP(CLK, M_EN, RST_M_DIV, M_DIV_END_OUT, M_OUT);

Z_GEN : FOR I IN 0 TO 6 GENERATE 
	    FF0 : IF(I = 0) GENERATE 
		        FFZ0 :FF PORT MAP(PDM_IN, REG_OUT(I), CLK, RST_ALL, LOAD);
				END GENERATE;
		FF1 : IF(I > 0) GENERATE		
	           FFZ1: FF PORT MAP(REG_OUT(I-1), REG_OUT(I), CLK, RST_ALL, LOAD);
			   END GENERATE;
        END GENERATE Z_GEN;

P0 : POLYPHASE_FIR GENERIC MAP(INITFILE => "POLYPHASE0.TXT") PORT MAP(CLK, RST_ALL, PDM_IN, M_DIV_END_IN, DAV0, POLY_VALID, P_OUT0);
P1 : POLYPHASE_FIR GENERIC MAP(INITFILE => "POLYPHASE1.TXT") PORT MAP(CLK, RST_ALL, REG_OUT(0), M_DIV_END_IN, DAV1, POLY_VALID, P_OUT1);
P2 : POLYPHASE_FIR GENERIC MAP(INITFILE => "POLYPHASE2.TXT") PORT MAP(CLK, RST_ALL, REG_OUT(1), M_DIV_END_IN, DAV2, POLY_VALID, P_OUT2);
P3 : POLYPHASE_FIR GENERIC MAP(INITFILE => "POLYPHASE3.TXT") PORT MAP(CLK, RST_ALL, REG_OUT(2), M_DIV_END_IN, DAV3, POLY_VALID, P_OUT3);
P4 : POLYPHASE_FIR GENERIC MAP(INITFILE => "POLYPHASE4.TXT") PORT MAP(CLK, RST_ALL, REG_OUT(3), M_DIV_END_IN, DAV4, POLY_VALID, P_OUT4);
P5 : POLYPHASE_FIR GENERIC MAP(INITFILE => "POLYPHASE5.TXT") PORT MAP(CLK, RST_ALL, REG_OUT(4), M_DIV_END_IN, DAV5, POLY_VALID, P_OUT5);
P6 : POLYPHASE_FIR GENERIC MAP(INITFILE => "POLYPHASE6.TXT") PORT MAP(CLK, RST_ALL, REG_OUT(5), M_DIV_END_IN, DAV6, POLY_VALID, P_OUT6);
P7 : POLYPHASE_FIR GENERIC MAP(INITFILE => "POLYPHASE7.TXT") PORT MAP(CLK, RST_ALL, REG_OUT(6), M_DIV_END_IN, DAV7, POLY_VALID, P_OUT7);


P_IN_MUX <= P_OUT7 & P_OUT6 & P_OUT5 & P_OUT4 & P_OUT3 & P_OUT2 & P_OUT1 & P_OUT0; --IN_MUX
DAV_OUT <= DAV7 & DAV6 & DAV5 & DAV4 & DAV3 & DAV2 & DAV1 & DAV0; 

MUX_SEL : N_COUNTER GENERIC MAP(N => 3, MODULE => 8) PORT MAP(CLK, EN_CNT_ADD, RST_ALL, CNT_END, CNT_OUT);

MUX: GENERICS_MUX GENERIC MAP(INPUTS => 8, SIZE => 28) PORT MAP(STD_LOGIC_VECTOR(P_IN_MUX), TO_INTEGER(CNT_OUT), P_OUT_MUX);

AS1 : ADD_SUB GENERIC MAP(N_AS => 28) PORT MAP(FILTER_OUT, SIGNED(P_OUT_MUX), AS_OUT, DAV_IN);

ACC_TOT : ACC GENERIC MAP(N_ACC => 28) PORT MAP(AS_OUT, FILTER_OUT, CLK, RST_ACC, EN_ACC);





END ARCHITECTURE;