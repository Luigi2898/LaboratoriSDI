LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY FIR IS
	GENERIC(INITFILE : STRING := "POLYPHASE.TXT");
	PORT(CLK         : IN STD_LOGIC; 
	     RST_FIR     : IN STD_LOGIC;
		 RST_CNT_FIR : IN STD_LOGIC;
	     EN_CNT_FIR  : IN STD_LOGIC; 		 
		 DOWNS_IN    : IN STD_LOGIC;
		 CNT_END_POLY: OUT STD_LOGIC; 	
		 OUT_MUX     : OUT STD_LOGIC_VECTOR(0 DOWNTO 0); 
		 PDM_AS      : IN STD_LOGIC;
		 EN_ACC      : IN STD_LOGIC;
		 RST_ACC     : IN STD_LOGIC;
		 LOAD_EN     : IN STD_LOGIC; 
		 SHIFT_EN    : IN STD_LOGIC; 
		 FIR_OUT     : BUFFER SIGNED(27 DOWNTO 0) 
	);
END ENTITY;


ARCHITECTURE BEH OF FIR IS

COMPONENT POLY_ROM IS
	GENERIC(INITFILE : STRING := "POLYPHASE.TXT";
	ADDR_N : INTEGER := 15; DATA_WIDTH : INTEGER := 20);
	PORT (CLK : IN STD_LOGIC;
		  ADDRESS : IN UNSIGNED(ADDR_N-1 DOWNTO 0);
		  DATAOUT : OUT SIGNED(DATA_WIDTH-1 DOWNTO 0)
	);
END COMPONENT; 
 
COMPONENT N_COUNTER IS
		GENERIC(N : INTEGER:= 6; MODULE : INTEGER := 42);
		PORT(CLK : IN STD_LOGIC;
			 EN  : IN STD_LOGIC;
			 RST : IN STD_LOGIC;
			 CNT_END : OUT STD_LOGIC;
			 CNT_OUT : BUFFER UNSIGNED(N-1 DOWNTO 0)		
		);
END COMPONENT;

COMPONENT SHIFTREGN IS
  GENERIC(
    N : INTEGER := 10
  );
  PORT (
    CLOCK    : IN STD_LOGIC;
    LOAD_EN  : IN STD_LOGIC;
    SHIFT_EN : IN STD_LOGIC;
    RSTN     : IN STD_LOGIC;    
	D_IN     : IN STD_LOGIC;
    D_OUT    : OUT STD_LOGIC;
	REG_OUT  : OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT GENERICS_MUX IS
	GENERIC(INPUTS : INTEGER := 15; SIZE: INTEGER := 1); --N INPUT, N BIT 
	PORT(INS : IN STD_LOGIC_VECTOR((INPUTS*SIZE)-1 DOWNTO 0);
		 SEL : IN INTEGER;
		 OUT_MUX : OUT STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0)
	);
END COMPONENT;

COMPONENT ACC IS 
	GENERIC(N_ACC : INTEGER := 14);
	PORT(ACC_IN : IN SIGNED(N_ACC-1 DOWNTO 0);
		 ACC_OUT : OUT SIGNED(N_ACC-1 DOWNTO 0);
		 CLK, RST, EN_ACC: IN STD_LOGIC	
	);
END COMPONENT;

COMPONENT ADD_SUB IS
	GENERIC(N_AS : INTEGER := 24);
	PORT(IN_AS_1, IN_AS_2 : IN SIGNED(N_AS-1 DOWNTO 0);
		 AS_OUT : OUT SIGNED(N_AS-1 DOWNTO 0);
		 PDM: IN STD_LOGIC
	);
END COMPONENT;

SIGNAL CNT_OUT_POLY: UNSIGNED(3 DOWNTO 0); --ADDRESS POLYPHASE
SIGNAL DOWNS_OUT: STD_LOGIC; --USCITA PDM SHIFT REG_OUT
SIGNAL SH_OUT : STD_LOGIC_VECTOR(12 DOWNTO 0); --SHIFT REG
SIGNAL POLY_OUT : SIGNED(27 DOWNTO 0);
SIGNAL AS_OUT: SIGNED(27 DOWNTO 0);

BEGIN 

P0 : POLY_ROM GENERIC MAP(INITFILE => INITFILE, ADDR_N => 4, DATA_WIDTH => 28) PORT MAP(CLK, CNT_OUT_POLY, POLY_OUT);

CNT: N_COUNTER GENERIC MAP(N => 4, MODULE => 13) PORT MAP(CLK, EN_CNT_FIR, RST_CNT_FIR, CNT_END_POLY, CNT_OUT_POLY);

SH : SHIFTREGN GENERIC MAP(N => 13) PORT MAP(CLK, LOAD_EN, SHIFT_EN, RST_FIR, DOWNS_IN, DOWNS_OUT, SH_OUT);

MUX : GENERICS_MUX GENERIC MAP(INPUTS => 13, SIZE => 1) PORT MAP(SH_OUT, TO_INTEGER(CNT_OUT_POLY), OUT_MUX);

AS : ADD_SUB GENERIC MAP(N_AS => 28) PORT MAP(FIR_OUT, POLY_OUT, AS_OUT, PDM_AS);

ACC1 : ACC GENERIC MAP(N_ACC => 28) PORT MAP(AS_OUT, FIR_OUT, CLK, RST_ACC, EN_ACC);








 

END ARCHITECTURE;