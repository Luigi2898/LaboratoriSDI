LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY CU_RX IS
	PORT(CLOCK         : IN STD_LOGIC;
         RST           : IN STD_LOGIC;		 
		 S_BIT         : IN STD_LOGIC;
		 DP_RST        : OUT STD_LOGIC;
		 RD            : OUT STD_LOGIC;
		 CNT1_EN       : OUT STD_LOGIC;
		 CNT1_END      : OUT STD_LOGIC;
		 CNT2_EN       : OUT STD_LOGIC;
		 CNT2_END      : OUT STD_LOGIC;
	     ENABLE_INPUT  : OUT STD_LOGIC;
		 ENABLE_OUTPUT : STD_LOGIC	
	);
END ENTITY;

ARCHITECTURE BEH OF CU_RX IS







END ARCHITECTURE;