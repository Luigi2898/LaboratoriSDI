LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;


ENTITY DP_FRONT_END IS
	PORT(CLK_10N : IN STD_LOGIC;
		 RST_CNT1 : IN STD_LOGIC;
		 RST_CNT2  : IN STD_LOGIC;
		 TC_HIGH : OUT STD_LOGIC;
		 TC_HIGH_NEG : OUT STD_LOGIC;
		 FF_IN : IN STD_LOGIC;
		 FF_OUT : OUT STD_LOGIC;
		 EN_FF1 : IN STD_LOGIC;
		 RST_FF1: IN STD_LOGIC;
		 FF_IN_NEG : IN STD_LOGIC;
		 FF_OUT_NEG : OUT STD_LOGIC;
		 EN_FF2  : IN STD_LOGIC;
		 RST_FF2 : IN STD_LOGIC
	);
END ENTITY;

ARCHITECTURE BEH OF DP_FRONT_END IS

COMPONENT RisingEdge_DFlipFlop_reset is
   port(
      Q : out std_logic;
      Clk :in std_logic;
      D :in  std_logic ;
      reset : in std_logic
   );
end COMPONENT;

COMPONENT N_COUNTER IS
		GENERIC(N : INTEGER:= 6; MODULE : INTEGER := 42);
		PORT(CLK : IN STD_LOGIC;
			 EN  : IN STD_LOGIC;
			 RST : IN STD_LOGIC;
			 CNT_END : OUT STD_LOGIC;
			 CNT_OUT : BUFFER UNSIGNED(N-1 DOWNTO 0)		
		);
END COMPONENT;

SIGNAL CNT_OUT1, CNT_OUT2 : UNSIGNED(5 DOWNTO 0);

BEGIN

TC1_HIGH : N_COUNTER GENERIC MAP(6, 47) PORT MAP(CLK_10N, EN_FF1, RST_CNT1, TC_HIGH, CNT_OUT1);

TC2_LOW : N_COUNTER GENERIC MAP(6, 47) PORT MAP(CLK_10N, EN_FF2, RST_CNT2, TC_HIGH_NEG, CNT_OUT2);

FF1 : RisingEdge_DFlipFlop_reset PORT MAP(FF_OUT, CLK_10N, FF_IN, RST_FF1);

FF2 : RisingEdge_DFlipFlop_reset PORT MAP(FF_OUT_NEG, CLK_10N, FF_IN_NEG, RST_FF2);


END ARCHITECTURE;


