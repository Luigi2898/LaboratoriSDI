LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

entity TB_POLYPHASE IS
END ENTITY;

ARCHITECTURE BEH OF TB_POLYPHASE IS

COMPONENT POLYPHASE_FIR IS
	GENERIC(INITFILE : STRING := "POLYPHASE.TXT");
	PORT(CLK        : IN STD_LOGIC;
	     RST        : IN STD_LOGIC;
	     DOWNS_IN   : IN STD_LOGIC;
	     M_DIV_END  : IN STD_LOGIC;
		 DAV        : OUT STD_LOGIC;
		 POLY_VALID : IN STD_LOGIC;
		 FIR_OUT    : BUFFER SIGNED(23 DOWNTO 0)
	);
END COMPONENT;


SIGNAL DOWNS_IN, M_DIV_END, POLY_VALID, DAV : STD_LOGIC;
SIGNAL FIR_OUT : SIGNED(23 DOWNTO 0);
SIGNAL RST, CLK: STD_LOGIC;

BEGIN

RST_PROCESS : PROCESS
BEGIN
	RST <= '0';
	WAIT FOR 5 NS;
	RST <= '1';
	wait for 20 sec;
END PROCESS;


clock : process
	begin
	
		clk <= '1';
		wait for 500 ns;
		clk <= '0';
		wait for 500 ns;
	
	end process;


P0 : POLYPHASE_FIR GENERIC MAP(INITFILE => "POLYPHASE0.TXT") PORT MAP(CLK, RST, DOWNS_IN, M_DIV_END, DAV, POLY_VALID, FIR_OUT);



END ARCHITECTURE;