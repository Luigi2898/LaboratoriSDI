library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity pippo is
  port (
  clock
  );
end entity;

architecture beh of pippo is

begin

end architecture;
